* /home/ahagen/scholarship/nucl_563/power_harvester/power_harvester.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue 18 Apr 2017 09:22:14 AM EDT

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
C2  2 11 4.7 uF		
C3  10 2 C		
C5  10 2 C		
C7  10 2 C		
C8  10 2 C		
L1  11 5 22 uH		
XU1  2 11 8 4 2 3 1 3 2 2 ? 2 2 10 10 5 2 BQ25504		
C4  2 10 4.7 uF		
C6  2 10 0.1 uF		
R3  1 3 R		
R4  3 2 R		
C1  4 2 0.01 uF		
R1  11 8 R		
R2  8 2 R		
D1  2 7 5 6 Diode_Bridge		

.end
